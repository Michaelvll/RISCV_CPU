`ifndef _IF
`define _IF

`include Defines
`include pc_reg

module IF (
    input wire clk,
    input wire rst,
    // input wire stall_s1_s2,
    // input wire pcsrc,
    // input wire jump_s4,
    // input wire baddr_s4,
    // input wire jaddr_s4,

    output reg [31:0]inst
);
    

endmodule





`endif