module cpu(
    input wire clk
);
// IF

// ID

// EX

// MEM

// WB

endmodule